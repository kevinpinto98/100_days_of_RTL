module tb_apb_slave();

endmodule