module tb_reg_file();


endmodule