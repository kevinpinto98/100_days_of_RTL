module tb_apb_master();


endmodule