module apb_master();


endmodule;