module tb_mem_interface();


endmodule