module apb_slave();


endmodule