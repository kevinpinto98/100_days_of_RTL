module d_ff();


endmodule
