module tb_rr_arbiter();


endmodule