module mem_interface();


endmodule