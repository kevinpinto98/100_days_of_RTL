module para_fifo();


endmodule