`timescale 1ns/100ps

module tb_dff();


endmodule
