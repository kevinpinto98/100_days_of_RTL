class day21;

function new();
//Nothing to do here
endfunction

function void print();
$display("Hi! This is day21 of the #100_day_RTL challenge");
endfunction

endclass