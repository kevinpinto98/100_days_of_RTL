module tb_para_fifo();


endmodule