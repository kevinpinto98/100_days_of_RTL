module day21_tb();

day21 Day21;

initial begin
    Day21 = new();
    Day21.print();
    $finish();
end


endmodule