module rr_arbiter();


endmodule